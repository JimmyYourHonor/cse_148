// sdram.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module sdram (
		input  wire        clk_clk,                              //                   clk.clk
		input  wire        d_cache_read_control_fixed_location,  //  d_cache_read_control.fixed_location
		input  wire [25:0] d_cache_read_control_read_base,       //                      .read_base
		input  wire [25:0] d_cache_read_control_read_length,     //                      .read_length
		input  wire        d_cache_read_control_go,              //                      .go
		output wire        d_cache_read_control_done,            //                      .done
		output wire        d_cache_read_control_early_done,      //                      .early_done
		input  wire        d_cache_read_user_read_buffer,        //     d_cache_read_user.read_buffer
		output wire [31:0] d_cache_read_user_buffer_output_data, //                      .buffer_output_data
		output wire        d_cache_read_user_data_available,     //                      .data_available
		input  wire        d_cache_write_control_fixed_location, // d_cache_write_control.fixed_location
		input  wire [25:0] d_cache_write_control_write_base,     //                      .write_base
		input  wire [25:0] d_cache_write_control_write_length,   //                      .write_length
		input  wire        d_cache_write_control_go,             //                      .go
		output wire        d_cache_write_control_done,           //                      .done
		input  wire        d_cache_write_user_write_buffer,      //    d_cache_write_user.write_buffer
		input  wire [31:0] d_cache_write_user_buffer_input_data, //                      .buffer_input_data
		output wire        d_cache_write_user_buffer_full,       //                      .buffer_full
		input  wire        i_cache_read_control_fixed_location,  //  i_cache_read_control.fixed_location
		input  wire [25:0] i_cache_read_control_read_base,       //                      .read_base
		input  wire [25:0] i_cache_read_control_read_length,     //                      .read_length
		input  wire        i_cache_read_control_go,              //                      .go
		output wire        i_cache_read_control_done,            //                      .done
		output wire        i_cache_read_control_early_done,      //                      .early_done
		input  wire        i_cache_read_user_read_buffer,        //     i_cache_read_user.read_buffer
		output wire [31:0] i_cache_read_user_buffer_output_data, //                      .buffer_output_data
		output wire        i_cache_read_user_data_available,     //                      .data_available
		output wire        mips_core_clk_clk,                    //         mips_core_clk.clk
		output wire        mips_core_rst_reset_n,                //         mips_core_rst.reset_n
		output wire        pll_0_locked_export,                  //          pll_0_locked.export
		input  wire        reset_reset_n,                        //                 reset.reset_n
		output wire        sdram_clk_clk,                        //             sdram_clk.clk
		output wire [12:0] sdram_controller_wire_addr,           // sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,             //                      .ba
		output wire        sdram_controller_wire_cas_n,          //                      .cas_n
		output wire        sdram_controller_wire_cke,            //                      .cke
		output wire        sdram_controller_wire_cs_n,           //                      .cs_n
		inout  wire [15:0] sdram_controller_wire_dq,             //                      .dq
		output wire [1:0]  sdram_controller_wire_dqm,            //                      .dqm
		output wire        sdram_controller_wire_ras_n,          //                      .ras_n
		output wire        sdram_controller_wire_we_n            //                      .we_n
	);

	wire  [31:0] d_cache_read_avalon_master_readdata;                 // mm_interconnect_0:d_cache_read_avalon_master_readdata -> d_cache_read:master_readdata
	wire         d_cache_read_avalon_master_waitrequest;              // mm_interconnect_0:d_cache_read_avalon_master_waitrequest -> d_cache_read:master_waitrequest
	wire  [25:0] d_cache_read_avalon_master_address;                  // d_cache_read:master_address -> mm_interconnect_0:d_cache_read_avalon_master_address
	wire         d_cache_read_avalon_master_read;                     // d_cache_read:master_read -> mm_interconnect_0:d_cache_read_avalon_master_read
	wire   [3:0] d_cache_read_avalon_master_byteenable;               // d_cache_read:master_byteenable -> mm_interconnect_0:d_cache_read_avalon_master_byteenable
	wire         d_cache_read_avalon_master_readdatavalid;            // mm_interconnect_0:d_cache_read_avalon_master_readdatavalid -> d_cache_read:master_readdatavalid
	wire         d_cache_write_avalon_master_waitrequest;             // mm_interconnect_0:d_cache_write_avalon_master_waitrequest -> d_cache_write:master_waitrequest
	wire  [25:0] d_cache_write_avalon_master_address;                 // d_cache_write:master_address -> mm_interconnect_0:d_cache_write_avalon_master_address
	wire   [3:0] d_cache_write_avalon_master_byteenable;              // d_cache_write:master_byteenable -> mm_interconnect_0:d_cache_write_avalon_master_byteenable
	wire         d_cache_write_avalon_master_write;                   // d_cache_write:master_write -> mm_interconnect_0:d_cache_write_avalon_master_write
	wire  [31:0] d_cache_write_avalon_master_writedata;               // d_cache_write:master_writedata -> mm_interconnect_0:d_cache_write_avalon_master_writedata
	wire  [31:0] i_cache_read_avalon_master_readdata;                 // mm_interconnect_0:i_cache_read_avalon_master_readdata -> i_cache_read:master_readdata
	wire         i_cache_read_avalon_master_waitrequest;              // mm_interconnect_0:i_cache_read_avalon_master_waitrequest -> i_cache_read:master_waitrequest
	wire  [25:0] i_cache_read_avalon_master_address;                  // i_cache_read:master_address -> mm_interconnect_0:i_cache_read_avalon_master_address
	wire         i_cache_read_avalon_master_read;                     // i_cache_read:master_read -> mm_interconnect_0:i_cache_read_avalon_master_read
	wire   [3:0] i_cache_read_avalon_master_byteenable;               // i_cache_read:master_byteenable -> mm_interconnect_0:i_cache_read_avalon_master_byteenable
	wire         i_cache_read_avalon_master_readdatavalid;            // mm_interconnect_0:i_cache_read_avalon_master_readdatavalid -> i_cache_read:master_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;    // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_readdata;      // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;   // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;       // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;          // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controller_s1_byteenable;    // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid; // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;         // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_writedata;     // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         rst_controller_reset_out_reset;                      // rst_controller:reset_out -> [d_cache_read:reset, d_cache_write:reset, i_cache_read:reset, mm_interconnect_0:d_cache_read_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_0:sdram_controller_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, sdram_controller:reset_n]

	custom_master #(
		.MASTER_DIRECTION    (0),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (26),
		.BURST_CAPABLE       (0),
		.MAXIMUM_BURST_COUNT (2),
		.BURST_COUNT_WIDTH   (2),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) d_cache_read (
		.clk                     (mips_core_clk_clk),                        //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),           // clock_reset_reset.reset
		.master_address          (d_cache_read_avalon_master_address),       //     avalon_master.address
		.master_read             (d_cache_read_avalon_master_read),          //                  .read
		.master_byteenable       (d_cache_read_avalon_master_byteenable),    //                  .byteenable
		.master_readdata         (d_cache_read_avalon_master_readdata),      //                  .readdata
		.master_readdatavalid    (d_cache_read_avalon_master_readdatavalid), //                  .readdatavalid
		.master_waitrequest      (d_cache_read_avalon_master_waitrequest),   //                  .waitrequest
		.control_fixed_location  (d_cache_read_control_fixed_location),      //           control.export
		.control_read_base       (d_cache_read_control_read_base),           //                  .export
		.control_read_length     (d_cache_read_control_read_length),         //                  .export
		.control_go              (d_cache_read_control_go),                  //                  .export
		.control_done            (d_cache_read_control_done),                //                  .export
		.control_early_done      (d_cache_read_control_early_done),          //                  .export
		.user_read_buffer        (d_cache_read_user_read_buffer),            //              user.export
		.user_buffer_output_data (d_cache_read_user_buffer_output_data),     //                  .export
		.user_data_available     (d_cache_read_user_data_available),         //                  .export
		.master_write            (),                                         //       (terminated)
		.master_writedata        (),                                         //       (terminated)
		.master_burstcount       (),                                         //       (terminated)
		.control_write_base      (26'b00000000000000000000000000),           //       (terminated)
		.control_write_length    (26'b00000000000000000000000000),           //       (terminated)
		.user_write_buffer       (1'b0),                                     //       (terminated)
		.user_buffer_input_data  (32'b00000000000000000000000000000000),     //       (terminated)
		.user_buffer_full        ()                                          //       (terminated)
	);

	custom_master #(
		.MASTER_DIRECTION    (1),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (26),
		.BURST_CAPABLE       (0),
		.MAXIMUM_BURST_COUNT (2),
		.BURST_COUNT_WIDTH   (2),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) d_cache_write (
		.clk                     (mips_core_clk_clk),                       //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),          // clock_reset_reset.reset
		.master_address          (d_cache_write_avalon_master_address),     //     avalon_master.address
		.master_write            (d_cache_write_avalon_master_write),       //                  .write
		.master_byteenable       (d_cache_write_avalon_master_byteenable),  //                  .byteenable
		.master_writedata        (d_cache_write_avalon_master_writedata),   //                  .writedata
		.master_waitrequest      (d_cache_write_avalon_master_waitrequest), //                  .waitrequest
		.control_fixed_location  (d_cache_write_control_fixed_location),    //           control.export
		.control_write_base      (d_cache_write_control_write_base),        //                  .export
		.control_write_length    (d_cache_write_control_write_length),      //                  .export
		.control_go              (d_cache_write_control_go),                //                  .export
		.control_done            (d_cache_write_control_done),              //                  .export
		.user_write_buffer       (d_cache_write_user_write_buffer),         //              user.export
		.user_buffer_input_data  (d_cache_write_user_buffer_input_data),    //                  .export
		.user_buffer_full        (d_cache_write_user_buffer_full),          //                  .export
		.master_read             (),                                        //       (terminated)
		.master_readdata         (32'b00000000000000000000000000000000),    //       (terminated)
		.master_readdatavalid    (1'b0),                                    //       (terminated)
		.master_burstcount       (),                                        //       (terminated)
		.control_read_base       (26'b00000000000000000000000000),          //       (terminated)
		.control_read_length     (26'b00000000000000000000000000),          //       (terminated)
		.control_early_done      (),                                        //       (terminated)
		.user_read_buffer        (1'b0),                                    //       (terminated)
		.user_buffer_output_data (),                                        //       (terminated)
		.user_data_available     ()                                         //       (terminated)
	);

	custom_master #(
		.MASTER_DIRECTION    (0),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (26),
		.BURST_CAPABLE       (0),
		.MAXIMUM_BURST_COUNT (2),
		.BURST_COUNT_WIDTH   (2),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) i_cache_read (
		.clk                     (mips_core_clk_clk),                        //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),           // clock_reset_reset.reset
		.master_address          (i_cache_read_avalon_master_address),       //     avalon_master.address
		.master_read             (i_cache_read_avalon_master_read),          //                  .read
		.master_byteenable       (i_cache_read_avalon_master_byteenable),    //                  .byteenable
		.master_readdata         (i_cache_read_avalon_master_readdata),      //                  .readdata
		.master_readdatavalid    (i_cache_read_avalon_master_readdatavalid), //                  .readdatavalid
		.master_waitrequest      (i_cache_read_avalon_master_waitrequest),   //                  .waitrequest
		.control_fixed_location  (i_cache_read_control_fixed_location),      //           control.export
		.control_read_base       (i_cache_read_control_read_base),           //                  .export
		.control_read_length     (i_cache_read_control_read_length),         //                  .export
		.control_go              (i_cache_read_control_go),                  //                  .export
		.control_done            (i_cache_read_control_done),                //                  .export
		.control_early_done      (i_cache_read_control_early_done),          //                  .export
		.user_read_buffer        (i_cache_read_user_read_buffer),            //              user.export
		.user_buffer_output_data (i_cache_read_user_buffer_output_data),     //                  .export
		.user_data_available     (i_cache_read_user_data_available),         //                  .export
		.master_write            (),                                         //       (terminated)
		.master_writedata        (),                                         //       (terminated)
		.master_burstcount       (),                                         //       (terminated)
		.control_write_base      (26'b00000000000000000000000000),           //       (terminated)
		.control_write_length    (26'b00000000000000000000000000),           //       (terminated)
		.user_write_buffer       (1'b0),                                     //       (terminated)
		.user_buffer_input_data  (32'b00000000000000000000000000000000),     //       (terminated)
		.user_buffer_full        ()                                          //       (terminated)
	);

	sdram_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (mips_core_clk_clk),   // outclk0.clk
		.outclk_1 (sdram_clk_clk),       // outclk1.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	sdram_sdram_controller sdram_controller (
		.clk            (mips_core_clk_clk),                                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	sdram_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                                          (mips_core_clk_clk),                                   //                                        pll_0_outclk0.clk
		.d_cache_read_clock_reset_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // d_cache_read_clock_reset_reset_reset_bridge_in_reset.reset
		.sdram_controller_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                      //         sdram_controller_reset_reset_bridge_in_reset.reset
		.d_cache_read_avalon_master_address                         (d_cache_read_avalon_master_address),                  //                           d_cache_read_avalon_master.address
		.d_cache_read_avalon_master_waitrequest                     (d_cache_read_avalon_master_waitrequest),              //                                                     .waitrequest
		.d_cache_read_avalon_master_byteenable                      (d_cache_read_avalon_master_byteenable),               //                                                     .byteenable
		.d_cache_read_avalon_master_read                            (d_cache_read_avalon_master_read),                     //                                                     .read
		.d_cache_read_avalon_master_readdata                        (d_cache_read_avalon_master_readdata),                 //                                                     .readdata
		.d_cache_read_avalon_master_readdatavalid                   (d_cache_read_avalon_master_readdatavalid),            //                                                     .readdatavalid
		.d_cache_write_avalon_master_address                        (d_cache_write_avalon_master_address),                 //                          d_cache_write_avalon_master.address
		.d_cache_write_avalon_master_waitrequest                    (d_cache_write_avalon_master_waitrequest),             //                                                     .waitrequest
		.d_cache_write_avalon_master_byteenable                     (d_cache_write_avalon_master_byteenable),              //                                                     .byteenable
		.d_cache_write_avalon_master_write                          (d_cache_write_avalon_master_write),                   //                                                     .write
		.d_cache_write_avalon_master_writedata                      (d_cache_write_avalon_master_writedata),               //                                                     .writedata
		.i_cache_read_avalon_master_address                         (i_cache_read_avalon_master_address),                  //                           i_cache_read_avalon_master.address
		.i_cache_read_avalon_master_waitrequest                     (i_cache_read_avalon_master_waitrequest),              //                                                     .waitrequest
		.i_cache_read_avalon_master_byteenable                      (i_cache_read_avalon_master_byteenable),               //                                                     .byteenable
		.i_cache_read_avalon_master_read                            (i_cache_read_avalon_master_read),                     //                                                     .read
		.i_cache_read_avalon_master_readdata                        (i_cache_read_avalon_master_readdata),                 //                                                     .readdata
		.i_cache_read_avalon_master_readdatavalid                   (i_cache_read_avalon_master_readdatavalid),            //                                                     .readdatavalid
		.sdram_controller_s1_address                                (mm_interconnect_0_sdram_controller_s1_address),       //                                  sdram_controller_s1.address
		.sdram_controller_s1_write                                  (mm_interconnect_0_sdram_controller_s1_write),         //                                                     .write
		.sdram_controller_s1_read                                   (mm_interconnect_0_sdram_controller_s1_read),          //                                                     .read
		.sdram_controller_s1_readdata                               (mm_interconnect_0_sdram_controller_s1_readdata),      //                                                     .readdata
		.sdram_controller_s1_writedata                              (mm_interconnect_0_sdram_controller_s1_writedata),     //                                                     .writedata
		.sdram_controller_s1_byteenable                             (mm_interconnect_0_sdram_controller_s1_byteenable),    //                                                     .byteenable
		.sdram_controller_s1_readdatavalid                          (mm_interconnect_0_sdram_controller_s1_readdatavalid), //                                                     .readdatavalid
		.sdram_controller_s1_waitrequest                            (mm_interconnect_0_sdram_controller_s1_waitrequest),   //                                                     .waitrequest
		.sdram_controller_s1_chipselect                             (mm_interconnect_0_sdram_controller_s1_chipselect)     //                                                     .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (mips_core_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	assign mips_core_rst_reset_n = ~rst_controller_reset_out_reset;

endmodule
